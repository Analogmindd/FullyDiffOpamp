** sch_path: /home/ubuntu/Desktop/FullyDiffOpamp/P_in_folded_cascode_RR_tb.sch
**.subckt P_in_folded_cascode_RR_tb
V2 GNDA 0 0
V5 VINP GNDA 0.7
V1 VINN GNDA 0.7
x1 net3 net4 VOUTN_BASE VOUTP_BASE VDDA GNDA VREF P_in_folded_cascode
V3 VDDA GNDA 1.8
V4 VREF GNDA 0.9
V6 net3 VINP AC 0.5
V7 net4 VINN AC -0.5
x2 VINP VINN VOUTN_PS VOUTP_PS net5 GNDA VREF P_in_folded_cascode
V8 net5 VDDA AC 1
x3 VINP VINN VOUTN_CM VOUTP_CM VDDA GNDA net1 P_in_folded_cascode
V9 net1 VREF AC 1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130B/libs.tech/ngspice/sky130.lib.spice ss



.control
save all
*op
ac dec 100 1 100T
setplot new
let frequency = ac.frequency
let T = ac.voutp_base-ac.voutn_base
let T_mag = db(T)
let T_ph  = cph(T)*180/pi

let T1 = ac.voutp_ps
let PSRR = T/T1
let PSRR_mag = db(PSRR)
let PSRR_ph  = cph(PSRR)*180/pi
let T1_mag = db(T1)
let T1_ph  = cph(T1)*180/pi
let T2 = (ac.voutp_cm-ac.voutn_cm)
let T2_mag = db(T2)
let T2_ph  = cph(T2)*180/pi
let CMRR = T/T2
let CMRR_mag = db(CMRR)
let CMRR_ph = cph(CMRR)*180/pi
plot T_mag T_ph xlog
plot T1_mag T1_ph xlog
plot PSRR_mag PSRR_ph xlog
plot CMRR_mag CMRR_ph xlog
write P_in_folded_cascode.raw
.endc

**** end user architecture code
**.ends

* expanding   symbol:  P_in_folded_cascode.sym # of pins=7
** sym_path: /home/ubuntu/Desktop/FullyDiffOpamp/P_in_folded_cascode.sym
** sch_path: /home/ubuntu/Desktop/FullyDiffOpamp/P_in_folded_cascode.sch
.subckt P_in_folded_cascode  VINP VINN VOUTN VOUTP VDDA GNDA VREF
*.ipin VINP
*.ipin VINN
*.opin VOUTN
*.opin VOUTP
*.ipin VDDA
*.ipin GNDA
*.ipin VREF
XM4 net1 VCMFB VDDA VDDA sky130_fd_pr__pfet_01v8_lvt L=0.7 W=11 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=60 m=60
XM5 net2 VCMFB VDDA VDDA sky130_fd_pr__pfet_01v8_lvt L=0.7 W=11 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=60 m=60
XM6 VOUTPF VB2 net1 VDDA sky130_fd_pr__pfet_01v8_lvt L=0.7 W=11.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
XM7 VOUTNF VB2 net2 VDDA sky130_fd_pr__pfet_01v8_lvt L=0.7 W=11.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
XM8 VOUTPF VB3 net3 GNDA sky130_fd_pr__nfet_01v8_lvt L=0.7 W=3.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=5 m=5
XM9 VOUTNF VB3 net4 GNDA sky130_fd_pr__nfet_01v8_lvt L=0.7 W=3.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=5 m=5
XM10 net3 VB4 net5 GNDA sky130_fd_pr__nfet_01v8_lvt L=0.7 W=2.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=9 m=9
XM11 net4 VB4 net5 GNDA sky130_fd_pr__nfet_01v8_lvt L=0.7 W=2.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=9 m=9
XM12 net6 VB1 VDDA VDDA sky130_fd_pr__pfet_01v8_lvt L=0.7 W=9.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=40 m=40
XM15 VB1 VB2 net6 VDDA sky130_fd_pr__pfet_01v8_lvt L=0.7 W=11.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
.save  v(vb1)
.save  v(net6)
R1 VB1 VB2 2.5k m=1
.save  v(vb2)
XM13 net7 VB4 net5 net5 sky130_fd_pr__nfet_01v8_lvt L=0.7 W=2.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=5 m=5
XM14 net8 VB4 net5 net5 sky130_fd_pr__nfet_01v8_lvt L=0.7 W=2.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=5 m=5
XM16 VB4 VB3 net7 net5 sky130_fd_pr__nfet_01v8_lvt L=0.7 W=3.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=5 m=5
XM17 VB2 VB3 net8 net5 sky130_fd_pr__nfet_01v8_lvt L=0.7 W=3.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=5 m=5
.save  v(net7)
.save  v(net8)
.save  v(vb4)
R2 VB3 VB4 2k m=1
I0 VDDA VB3 200u
XM18 VOUTN VOUTPF net5 net5 sky130_fd_pr__nfet_01v8_lvt L=0.7 W=14.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=21 m=21
XM19 VOUTN net9 VDDA VDDA sky130_fd_pr__pfet_01v8_lvt L=0.7 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=66 m=66
XM20 VOUTP VOUTNF net5 net5 sky130_fd_pr__nfet_01v8_lvt L=0.7 W=14.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=21 m=21
XM21 VOUTP net9 VDDA VDDA sky130_fd_pr__pfet_01v8_lvt L=0.7 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=66 m=66
R5 net10 VOUTPF 100 m=1
R6 net11 VOUTNF 100 m=1
C1 VOUTN net10 1.1p m=1
C2 VOUTP net11 1.1p m=1
.save  v(net1)
.save  v(net2)
.save  v(voutpf)
.save  v(voutnf)
.save  v(net3)
.save  v(net4)
.save  v(voutn)
.save  v(voutp)
.save  v(vb3)
XM1 net12 VB1 VDDA VDDA sky130_fd_pr__pfet_01v8_lvt L=0.7 W=9.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=58 m=58
XM2 net3 VINN net12 VDDA sky130_fd_pr__pfet_01v8_lvt L=0.7 W=10.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=20 m=20
XM3 net12 VINP net4 VDDA sky130_fd_pr__pfet_01v8_lvt L=0.7 W=10.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=20 m=20
R3 net9 VOUTN 100Meg m=1
R4 VOUTP net9 100Meg m=1
XM22 net13 VB4 net5 net5 sky130_fd_pr__nfet_01v8_lvt L=0.7 W=2.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM23 net14 VB4 net5 net5 sky130_fd_pr__nfet_01v8_lvt L=0.7 W=2.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM24 VCMFB VREF net13 GNDA sky130_fd_pr__nfet_01v8_lvt L=0.7 W=14.1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM25 VCMFB VREF net14 GNDA sky130_fd_pr__nfet_01v8_lvt L=0.7 W=14.1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM26 net15 VOUTPF net13 GNDA sky130_fd_pr__nfet_01v8_lvt L=0.7 W=14.1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM27 net15 VOUTNF net14 GNDA sky130_fd_pr__nfet_01v8_lvt L=0.7 W=14.1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM28 VCMFB VCMFB VDDA VDDA sky130_fd_pr__pfet_01v8_lvt L=0.7 W=11 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
XM29 net15 net15 VDDA VDDA sky130_fd_pr__pfet_01v8_lvt L=0.7 W=11 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
.save  v(net13)
.save  v(net14)
.save  v(vcmfb)
.save  v(net15)
.save  v(net9)
C7 VOUTP GNDA 5p m=1
C8 VOUTN GNDA 5p m=1
Vmeas net5 GNDA 0
.save  i(vmeas)
.ends

.end
